module connection(
	input wire in_1,
	output wire out_1
);
assign out_1=in_1;
endmodule
